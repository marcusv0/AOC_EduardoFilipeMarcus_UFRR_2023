-----------------------------------------------------------
-- COMPONENTE: MEMÓRIA ROM
-- DESCRIÇÃO: 
--     RESPONSÁVEL POR ARMAZENAR O PROGRAMA A SER EXECUTADO
--     UTILIZANDO DA SEGUINTE SINTAXE:
--     TIPO R:
--	   | OPCODE "XXXX" | RS "XX" | RT "XX" |
--     TIPO I:
--         | OPCODE "XXXX" | RS "XX" | VALOR "XX |
--     TIPO J:
--	   | OPCODE "XXXX" | ENDEREÇO "XXXX" |
--     ESSAS INSTRUÇÕES DO PROGRAMA SÃO ARMAZENADAS NOS 256
--     BYTES DE MEMÓRIA DISPONÍVEIS
-----------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ROM IS
    PORT(
        CLOCK : IN STD_LOGIC;
        A     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        S     : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE BEHAVIOR OF ROM IS
    TYPE MEM_T IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
    CONSTANT MEM : MEM_T := (
-- PARA EXECUTAR OS TESTES É SÓ TIRAR O COMENTÁRIO
	
-- TESTE DE SUB E SUBI
--		0 => "0000000000010011", -- ADDI S0 3
--		1 => "0000000000010101", -- ADDI S1 1
--		2 => "0000000001100001", -- SUBI S0 1
--		3 => "0000000001000001", -- SUB S0 S1

-- TESTE DE ADD E ADDI
--		0 => "0000000000010011", -- ADDI S0 3
--		1 => "0000000000010111", -- ADDI S1 3
--		2 => "0000000000000001", -- ADD S0 S1
		
-- TESTE BEQ
--		0 => "0000000001100010", -- LI S0 2
--		1 => "0000000001100110", -- LI S1 2
--		2 => "0000000100000001", -- IF S0 == S1
--		3 => "0000000001110101", -- BEQ S0 == S1 JUMP 0101
--		4 => "0000000000010001", -- ADDI S0 1
--		5 => "0000000000010010", -- ADDI S0 2

-- TESTE LI
--		0 => "0000000001100010", -- LI S0 2
--		1 => "0000000000000001", -- ADDI S0 1

		
-- TESTE FIBONACCI
--		0 => "0000000000010000", -- ADDI S0 0
--		1 => "0000000001010000", -- SW S0
--		2 => "0000000000010001", -- ADDI S0 1
--		3 => "0000000000010101", -- ADDI S1 1
--		4 => "0000000001001100", -- LW S3 00
--		5 => "0000000000101101", -- ADD S3 S1
--		6 => "0000000000000100", -- ADD S1 S0
--		7 => "0000000001000000", -- LW S0 00
--		8 => "0000000000000011", -- ADD S0 S3
--		9 => "0000000001010100", -- J 0100

      OTHERS => "0000000001111111"
    );
BEGIN
    PROCESS(CLOCK, A)
    BEGIN
        S <= MEM(CONV_INTEGER(UNSIGNED(A(15 DOWNTO 8))));
    END PROCESS;
END;
