-----------------------------------------------------------
-- COMPONENTE: MEMÓRIA ROM
-- DESCRIÇÃO: 
--     RESPONSÁVEL POR ARMAZENAR O PROGRAMA A SER EXECUTADO
--     0001 000000 00011
-----------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY ROM IS
    PORT(
        CLOCK : IN STD_LOGIC;
        A     : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        S     : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE BEHAVIOR OF ROM IS
    TYPE MEM_T IS ARRAY (0 TO 255) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
    CONSTANT MEM : MEM_T := (
-- PARA EXECUTAR RETIRE O COMENTÁRIO

---- TESTE DE ADDI, SUB E SUBI
--		0 => "0001000000000011", -- ADDI S0 3
--		1 => "0001000001000001", -- ADDI S1 1
--		2 => "0011000000000001", -- SUBI S0 1
--		3 => "0010000000000001", -- SUB S0 S1

---- TESTE DE ADD E ADDI
--		0 => "0001000000000011", -- ADDI S0 3
--		1 => "0001000001000011", -- ADDI S1 3
--		2 => "0000000000000001", -- ADD S0 S1
		
---- TESTE BEQ
--		0 => "0110000000000010", -- LI S0 2
--		1 => "0110000001000010", -- LI S1 2
--		2 => "1000000000000001", -- IF S0 == S1
--		3 => "0111000000000101", -- BEQ S0 == S1 JUMP 
--		4 => "0001000000000001", -- ADDI S0 1
--		5 => "0001000000000010", -- ADDI S0 2

-- -- TESTE LI
--		0 => "0110000000000010", -- LI S0 2
--		1 => "0001000000000001", -- ADDI S0 1

		
-- TESTE FIBONACCI
		0 => "0001000000000000", -- ADDI S0 0
		1 => "0101000000000000", -- SW S0
		2 => "0001000000000001", -- ADDI S0 1
		3 => "0001000001000001", -- ADDI S1 1
		4 => "0100000010000000", -- LW S2 0
		5 => "0000000010000001", -- ADD S2 S1
		6 => "0000000000000000", -- ADD S1 S0
		7 => "0100000001000000", -- LW S0 00
		8 => "0000000000000010", -- ADD S0 S2
		9 => "1001000001010100", -- J 0100

      OTHERS => "0000000001111111"
    );
BEGIN
    PROCESS(CLOCK, A)
    BEGIN
        S <= MEM(CONV_INTEGER(UNSIGNED(A)));
    END PROCESS;
END;
